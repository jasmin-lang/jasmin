(** This module is meant as the minimal dependency of extracted code. *)
From compiler Require compiler.
From lang Require psem_defs.
From armv7 Require arm_params.
From x86 Require x86_params.
From riscv Require riscv_params.
From arch Require sem_params_of_arch_extra.
From compiler Require wint_int.

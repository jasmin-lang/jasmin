(** This module is meant as the minimal dependency of extracted code. *)
Require compiler.
Require psem_defs.
Require arm_params.
Require x86_params.
Require riscv_params.
Require sem_params_of_arch_extra.
Require safety_cond.
Require contracts_asserts.
Require remove_is_var_init.
Require extra_vars_call.

